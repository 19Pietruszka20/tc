module test ;
initial begin
$display ( " Hello World ! " );
end
endmodule